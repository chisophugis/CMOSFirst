*** SPICE deck for cell inverter_sim{lay} from library tutorial_4
*** Created on Sun Feb 15, 2015 15:26:46
*** Last revised on Sun Feb 15, 2015 15:36:08
*** Written on Tue Feb 17, 2015 22:15:27 by Electric VLSI Design System,
*** version 9.05
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT tutorial_4__inv_20_10 FROM CELL inv_20_10{lay}
.SUBCKT tutorial_4__inv_20_10 gnd in out vdd
Mnmos@0 out in gnd gnd myNMOS L=0.2U W=6U AS=14.4P AD=8.1P PS=24.6U PD=12.6U
Mpmos@0 out in vdd vdd myPMOS L=0.2U W=12U AS=19.8P AD=8.1P PS=30.6U PD=12.6U
.ENDS tutorial_4__inv_20_10

*** TOP LEVEL CELL: inverter_sim{lay}
Xinv_20_1@0 gnd inwire outwire vdd tutorial_4__inv_20_10

Xinv_20_1@1 gnd outwire outwire2 vdd tutorial_4__inv_20_10

Xinv_20_1@2 gnd outwire2 outwire3 vdd tutorial_4__inv_20_10
Xinv_20_1@3 gnd outwire3 outwire4 vdd tutorial_4__inv_20_10
Xinv_20_1@4 gnd outwire4 inwire vdd tutorial_4__inv_20_10

* Xinv_20_1@3 gnd outwire3 inwire vdd tutorial_4__inv_20_10

* Spice Code nodes in cell cell 'inverter_sim{lay}'
vdd vdd 0 DC 5
*vin vin 0 PULSE(0 5 100p)
*r1 vin inwire 10k


*vin inwire 0 PULSE(0 5 100p 50p 50p 300p)
.ic V(inwire)=0
*.dc vin 0 5 1m
.tran 10000p uic
.include C5_models.txt
.END
